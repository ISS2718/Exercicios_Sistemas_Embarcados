-- ###################################################################################################
-- # << ISS2718 - Top Level File for Matrix Multiplication Accelerator >>                            #
-- # *********************************************************************************************** #
-- # NOTE: This is a custom subsystem for accelerating matrix multiplication,                        #
-- # through a scalar product hardware accelerator.                                                  #
-- #                                                                                                 #
-- #       This code is a modification of the NEORV32 RISC-V Processor,                              #
-- #       available at https://github.com/stnolting/neorv32                                         #
-- #       Modified by Daniel Contente, Hugo Nakamura, Isaac Soares, Mateus Messias                  #
-- # *********************************************************************************************** #
-- # BSD 3-Clause License                                                                            #
-- #                                                                                                 #
-- # Hardware matrix accelerator,                                                                    #
-- # https://github.com/ISS2718/Sistemas_Embarcados/Coprocessador                                    #
-- #                                                                                                 #
-- # Copyright (c) 2024, Daniel Contente, Hugo Nakamura, Isaac Soares, Mateus Messias. All rights    #
-- # reserved.                                                                                       #
-- #                                                                                                 #
-- # Redistribution and use in source and binary forms, with or without modification, are            #
-- # permitted provided that the following conditions are met:                                       #
-- #                                                                                                 #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of          #
-- #    conditions and the following disclaimer.                                                     #
-- #                                                                                                 #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of       #
-- #    conditions and the following disclaimer in the documentation and/or other materials          #
-- #    provided with the distribution.                                                              #
-- #                                                                                                 #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to    #
-- #    endorse or promote products derived from this software without specific prior written        #
-- #    permission.                                                                                  #
-- #                                                                                                 #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS     #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY #
-- # AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER     #
-- # OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR          #
-- # CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR        #
-- # SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY    #
-- # THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE       #
-- # OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE        #
-- # POSSIBILITY OF SUCH DAMAGE.                                                                     #
-- ###################################################################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library neorv32;
use neorv32.neorv32_package.all;

entity neorv32_matrix_accelerator is
  generic (
    -- adapt these for your setup --
    CLOCK_FREQUENCY   : natural := 50000000;  -- clock frequency of clk_i in Hz
    MEM_INT_IMEM_SIZE : natural := 64*1024;   -- size of processor-internal instruction memory in bytes
    MEM_INT_DMEM_SIZE : natural := 512*1024   -- size of processor-internal data memory in bytes
  );
  port (
    -- Global control --
    clk_i       : in  std_ulogic; -- global clock, rising edge
    rstn_i      : in  std_ulogic; -- global reset, low-active, async
    -- GPIO --
    gpio_o      : out std_ulogic_vector(7 downto 0); -- parallel output
    -- UART0 --
    uart0_txd_o : out std_ulogic; -- UART0 send data
    uart0_rxd_i : in  std_ulogic  -- UART0 receive data
  );
end entity;

architecture neorv32_test_setup_bootloader_rtl of neorv32_matrix_accelerator is

  signal con_gpio_o : std_ulogic_vector(63 downto 0);

begin

  -- The Core Of The Problem ----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  neorv32_top_inst: neorv32_top
  generic map (
    -- General --
    CLOCK_FREQUENCY              => CLOCK_FREQUENCY,   -- clock frequency of clk_i in Hz
    INT_BOOTLOADER_EN            => true,              -- boot configuration: true = boot explicit bootloader; false = boot from int/ext (I)MEM
    -- RISC-V CPU Extensions --
    CPU_EXTENSION_RISCV_C        => true,              -- implement compressed extension?
    CPU_EXTENSION_RISCV_M        => true,              -- implement mul/div extension?
    CPU_EXTENSION_RISCV_Zicntr   => true,              -- implement base counters?
    -- Internal Instruction memory --
    MEM_INT_IMEM_EN              => true,              -- implement processor-internal instruction memory
    MEM_INT_IMEM_SIZE            => MEM_INT_IMEM_SIZE, -- size of processor-internal instruction memory in bytes
    -- Internal Data memory --
    MEM_INT_DMEM_EN              => true,              -- implement processor-internal data memory
    MEM_INT_DMEM_SIZE            => MEM_INT_DMEM_SIZE, -- size of processor-internal data memory in bytes
    -- Processor peripherals --
    IO_GPIO_NUM                  => 8,                 -- number of GPIO input/output pairs (0..64)
    IO_MTIME_EN                  => true,              -- implement machine system timer (MTIME)?
    IO_UART0_EN                  => true,              -- implement primary universal asynchronous receiver/transmitter (UART0)?

    -- Custom Functions Subsystem --
    IO_CFS_EN                    => true,              -- implement custom functions subsystem (CFS)?
    IO_CFS_IN_SIZE               => 32,                -- size of CFS input conduit in bits
    IO_CFS_OUT_SIZE              => 32                -- size of CFS output conduit in bits
 )
  port map (
    -- Global control --
    clk_i       => clk_i,       -- global clock, rising edge
    rstn_i      => rstn_i,      -- global reset, low-active, async
    -- GPIO (available if IO_GPIO_EN = true) --
    gpio_o      => con_gpio_o,  -- parallel output
    -- primary UART0 (available if IO_GPIO_NUM > 0) --
    uart0_txd_o => uart0_txd_o, -- UART0 send data
    uart0_rxd_i => uart0_rxd_i  -- UART0 receive data
  );

  -- GPIO output --
  gpio_o <= con_gpio_o(7 downto 0);


end architecture;
